LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ABS_FSM_BLOCK IS
	GENERIC(TAU : TIME := 30 ps);
	PORT(
		CLK,RES : IN STD_LOGIC;
		FBP, RBP : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		FRS,FLS,RRS,RLS : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		SPD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		ABS_STATUS_F : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		ABS_STATUS_R : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END ENTITY ABS_FSM_BLOCK;

ARCHITECTURE RTL OF ABS_FSM_BLOCK IS
TYPE STATUS_F IS (IDLE,FBMS,FFLS,FRWSS,FLWSS,ERRS);
TYPE STATUS_R IS (IDLE,RBMS,FRLS,RRWSS,RLWSS,ERRS);
SIGNAL STATE_NOW_REAR, STATE_NEXT_REAR : STATUS_R;
SIGNAL STATE_NOW_FRONT, STATE_NEXT_FRONT : STATUS_F;
SIGNAL FULL_LOCK : STD_LOGIC := '0';
BEGIN
 PROCESS(CLK,RES)
  BEGIN
	IF(RES='1')THEN
		FULL_LOCK<='0';
		STATE_NOW_REAR<=IDLE;
		STATE_NOW_FRONT<=IDLE;
	ELSIF(RISING_EDGE(CLK))THEN 
		STATE_NOW_REAR<=STATE_NEXT_REAR;
		STATE_NOW_FRONT<=STATE_NEXT_FRONT;
	END IF;
 END PROCESS;
 
 PROCESS(STATE_NOW_FRONT,FBP)
  CONSTANT BRAKE_THRESHOLD : STD_LOGIC_VECTOR(2 DOWNTO 0) := "110";
  CONSTANT MOVING : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
  CONSTANT FULL_STOP : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
  CONSTANT SPEED_THRESHOLD : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
  CONSTANT SPINNING_TOLERANCE : REAL := 1.8;
  BEGIN
  	CASE STATE_NOW_FRONT IS
		WHEN IDLE =>
			IF(TO_INTEGER(UNSIGNED(SPD))>TO_INTEGER(UNSIGNED(MOVING)))THEN 
				STATE_NEXT_FRONT<=FBMS;
			ELSIF(STATE_NEXT_FRONT=FFLS) THEN
				STATE_NEXT_FRONT<=ERRS;
			END IF;
		WHEN FBMS =>
			IF(TO_INTEGER(UNSIGNED(FBP))>TO_INTEGER(UNSIGNED(BRAKE_THRESHOLD))) THEN
				STATE_NEXT_FRONT<=FFLS;
			ELSIF(((REAL(TO_INTEGER(UNSIGNED(FRS)))/(SPINNING_TOLERANCE))>REAL(TO_INTEGER(UNSIGNED(FLS)))) AND (TO_INTEGER(UNSIGNED(SPD))>(TO_INTEGER(UNSIGNED(SPEED_THRESHOLD))))) THEN
				STATE_NEXT_FRONT<=FRWSS;
			ELSIF(((REAL(TO_INTEGER(UNSIGNED(FLS)))/(SPINNING_TOLERANCE))>REAL(TO_INTEGER(UNSIGNED(FRS)))) AND (TO_INTEGER(UNSIGNED(SPD))>(TO_INTEGER(UNSIGNED(SPEED_THRESHOLD))))) THEN
				STATE_NEXT_FRONT<=FLWSS;
			ELSIF(TO_INTEGER(UNSIGNED(SPD))=(TO_INTEGER(UNSIGNED(FULL_STOP)))) THEN
				STATE_NEXT_FRONT<=IDLE;
			END IF;
		WHEN FFLS =>
			IF(TO_INTEGER(UNSIGNED(FBP))<TO_INTEGER(UNSIGNED(BRAKE_THRESHOLD))) THEN
				STATE_NEXT_FRONT<=FBMS;
			ELSIF(TO_INTEGER(UNSIGNED(SPD))=(TO_INTEGER(UNSIGNED(FULL_STOP)))) THEN
				STATE_NEXT_FRONT<=IDLE;
			END IF;
		WHEN FRWSS =>
			IF(((REAL(TO_INTEGER(UNSIGNED(FRS)))/(SPINNING_TOLERANCE))<REAL(TO_INTEGER(UNSIGNED(FLS)))) OR (TO_INTEGER(UNSIGNED(SPD))<(TO_INTEGER(UNSIGNED(SPEED_THRESHOLD))))) THEN
				STATE_NEXT_FRONT<=FBMS;
			ELSIF(TO_INTEGER(UNSIGNED(SPD))=(TO_INTEGER(UNSIGNED(FULL_STOP)))) THEN
				STATE_NEXT_FRONT<=IDLE;
			END IF;
		WHEN FLWSS =>
			IF(((REAL(TO_INTEGER(UNSIGNED(FLS)))/(SPINNING_TOLERANCE))<REAL(TO_INTEGER(UNSIGNED(FRS)))) OR (TO_INTEGER(UNSIGNED(SPD))<(TO_INTEGER(UNSIGNED(SPEED_THRESHOLD))))) THEN
				STATE_NEXT_FRONT<=FBMS;
			ELSIF(TO_INTEGER(UNSIGNED(SPD))=(TO_INTEGER(UNSIGNED(FULL_STOP)))) THEN
				STATE_NEXT_FRONT<=IDLE;
			END IF;
		WHEN OTHERS =>
			NULL;
	END CASE;
 END PROCESS;

 PROCESS(STATE_NOW_REAR,RBP)
  CONSTANT BRAKE_THRESHOLD : STD_LOGIC_VECTOR(2 DOWNTO 0) := "110";
  CONSTANT MOVING : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
  CONSTANT FULL_STOP : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
  CONSTANT SPEED_THRESHOLD : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
  CONSTANT SPINNING_TOLERANCE : REAL := 1.8;
  BEGIN
  	CASE STATE_NOW_REAR IS
		WHEN IDLE =>
			IF(TO_INTEGER(UNSIGNED(SPD))>TO_INTEGER(UNSIGNED(MOVING)))THEN 
				STATE_NEXT_REAR<=RBMS;
			ELSIF(STATE_NEXT_REAR=FRLS) THEN 
  				STATE_NEXT_REAR<=ERRS;
			END IF;
		WHEN RBMS =>
			IF(TO_INTEGER(UNSIGNED(RBP))>TO_INTEGER(UNSIGNED(BRAKE_THRESHOLD))) THEN
				STATE_NEXT_REAR<=FRLS;
			ELSIF(((REAL(TO_INTEGER(UNSIGNED(RRS)))/(SPINNING_TOLERANCE))>REAL(TO_INTEGER(UNSIGNED(RLS)))) AND (TO_INTEGER(UNSIGNED(SPD))>(TO_INTEGER(UNSIGNED(SPEED_THRESHOLD))))) THEN
				STATE_NEXT_REAR<=RRWSS;
			ELSIF(((REAL(TO_INTEGER(UNSIGNED(RLS)))/(SPINNING_TOLERANCE))>REAL(TO_INTEGER(UNSIGNED(FRS)))) AND (TO_INTEGER(UNSIGNED(SPD))>(TO_INTEGER(UNSIGNED(SPEED_THRESHOLD))))) THEN
				STATE_NEXT_REAR<=RLWSS;
			ELSIF(TO_INTEGER(UNSIGNED(SPD))=(TO_INTEGER(UNSIGNED(FULL_STOP)))) THEN
				STATE_NEXT_REAR<=IDLE;
			END IF;
		WHEN FRLS =>
			IF(TO_INTEGER(UNSIGNED(RBP))<TO_INTEGER(UNSIGNED(BRAKE_THRESHOLD))) THEN
				STATE_NEXT_REAR<=RBMS;
			ELSIF(TO_INTEGER(UNSIGNED(SPD))=(TO_INTEGER(UNSIGNED(FULL_STOP)))) THEN
				STATE_NEXT_REAR<=IDLE;
			END IF;
		WHEN RRWSS =>
			IF(((REAL(TO_INTEGER(UNSIGNED(RRS)))/(SPINNING_TOLERANCE))<REAL(TO_INTEGER(UNSIGNED(RLS)))) OR (TO_INTEGER(UNSIGNED(SPD))<(TO_INTEGER(UNSIGNED(SPEED_THRESHOLD))))) THEN
				STATE_NEXT_REAR<=RBMS;
			ELSIF(TO_INTEGER(UNSIGNED(SPD))=(TO_INTEGER(UNSIGNED(FULL_STOP)))) THEN
				STATE_NEXT_REAR<=IDLE;
			END IF;
		WHEN RLWSS =>
			IF(((REAL(TO_INTEGER(UNSIGNED(RLS)))/(SPINNING_TOLERANCE))<REAL(TO_INTEGER(UNSIGNED(RRS)))) OR (TO_INTEGER(UNSIGNED(SPD))<(TO_INTEGER(UNSIGNED(SPEED_THRESHOLD))))) THEN
				STATE_NEXT_REAR<=RBMS;
			ELSIF(TO_INTEGER(UNSIGNED(SPD))=(TO_INTEGER(UNSIGNED(FULL_STOP)))) THEN
				STATE_NEXT_REAR<=IDLE;
			END IF;
		WHEN OTHERS =>
			NULL;
	END CASE;
 END PROCESS;
 -- psl endpoints to evaluate states useful for assertions
 --psl endpoint E_FFLS_FBMS is {STATE_NOW_FRONT = FFLS; STATE_NOW_FRONT = FBMS}@CLK'active;
 --psl endpoint E_FRLS_RBMS is {STATE_NOW_REAR = FRLS; STATE_NOW_REAR = RBMS}@CLK'active;
 --psl endpoint E_ERRS_R is {STATE_NOW_REAR = ERRS}@CLK'active;
 --psl endpoint E_ERRS_F is {STATE_NOW_FRONT = ERRS}@CLK'active;

 -- Determining the full lock state
 PROCESS(STATE_NOW_REAR,STATE_NOW_FRONT)
 BEGIN
	IF (STATE_NOW_REAR=FRLS AND STATE_NOW_FRONT=FFLS) THEN
		FULL_LOCK<='1';
	ELSE FULL_LOCK <= '0';
	END IF;
 END PROCESS;
 -- Output process 
 PROCESS(STATE_NOW_REAR,STATE_NOW_FRONT)
  BEGIN
  	
  	IF (FULL_LOCK='1') THEN
  		ABS_STATUS_F<="1111" AFTER TAU;
  		ABS_STATUS_R<="1111" AFTER TAU;
	ELSE
		CASE STATE_NOW_FRONT IS
			WHEN FBMS =>
				ABS_STATUS_F<="0001" AFTER TAU;
			WHEN FFLS =>
				ABS_STATUS_F<="0010" AFTER TAU;
			WHEN FRWSS =>
				ABS_STATUS_F<="0011" AFTER TAU;
			WHEN FLWSS =>
				ABS_STATUS_F<="0100" AFTER TAU;
			WHEN ERRS =>
				ABS_STATUS_F<="0101" AFTER TAU;
			WHEN IDLE =>
				ABS_STATUS_F<="0000" AFTER TAU;
		END CASE;
		CASE STATE_NOW_REAR IS
			WHEN RBMS =>
				ABS_STATUS_R<="1110" AFTER TAU;
			WHEN FRLS =>
				ABS_STATUS_R<="1101" AFTER TAU;
			WHEN RRWSS =>
				ABS_STATUS_R<="1100" AFTER TAU;
			WHEN RLWSS =>
				ABS_STATUS_R<="1011" AFTER TAU;
			WHEN ERRS =>
				ABS_STATUS_R<="0101" AFTER TAU;
			WHEN IDLE =>
				ABS_STATUS_R<="0000" AFTER TAU;
		END CASE;
	END IF;
 END PROCESS;

 --psl default clock is rising_edge(CLK);
 --psl property anti_full_lock is always (FULL_LOCK -> next![3](not(FULL_LOCK)));
 --psl property anti_front_lock is always (STATE_NOW_FRONT = FFLS) -> next[3](STATE_NOW_FRONT=FBMS);
 --psl property anti_rear_lock is always ((STATE_NOW_REAR=FRLS) -> next[3](STATE_NOW_REAR=RBMS));
 --psl property anti_errs_r is always ((STATE_NOW_REAR=ERRS) -> next![3](not(STATE_NOW_REAR=ERRS)));
 --psl property anti_errs_f is always ((STATE_NOW_FRONT=ERRS) -> next![3](not(STATE_NOW_FRONT=ERRS)));

 --psl assert anti_full_lock;
 --psl assert anti_front_lock;
 --psl assert anti_rear_lock;
 --psl assert anti_errs_f;
END ARCHITECTURE RTL;
			
